// CN1 -  schelet lab02
// structural
module modul01(
  output out,
  input in
  );

  not(out, in);

endmodule