module ex1(
    output  AN0,
    output  AN1,
    output  AN2,
    output  AN3,
    output  CA,
    output  CB,
    output  CC,
    output  CD,
    output  CE,
    output  CF,
    output  CG,
    output  DP
    );

    // TODO
	 assign AN0 = 0;
	 assign AN1 = 0;
	 assign AN2 = 0;
	 assign AN3 = 0;
	 assign CA = 0;
	 assign CB = 0;
	 assign CG = 1;
	 assign CC = 0;
	 assign CD = 0;
	 assign CE = 0;
	 assign CF = 0;
	 assign DP = 1;
	 
endmodule
